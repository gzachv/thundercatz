/****************************************************************
 Module to implement the circular queue opperating at 24.424kHz.
 Authors : ThunderCatz 		HDL : System Verilog		 
 Student ID: 903 015 5247	
 Date : 11/13/2015 							
****************************************************************/ 

////////// Variable Declaration for interface ///////////////////

////////// Intermediate wire Declarations ///////////////////////
